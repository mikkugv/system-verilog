module tb;
    integer_example uut();
    initial begin
        #50;
        $finish;
    end
endmodule
